`define simulation