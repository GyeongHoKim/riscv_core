//`define simulation
// do not define when you work on fpga, do define when you simulate